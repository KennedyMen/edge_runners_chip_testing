module test (
    input [7:0] in,
    out,
    input clk,
    rst,
    input en
);


endmodule
