module Mensah (
  ports
   heloo
);
  
