module sqrt_22b (
    input  logic [21:0] value,     
    output logic [10:0] sqrt    
);
    

    const logic [10:0] sqrt_below_1024 [0:1023] = '{
        0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32
    };

    const logic [10:0] sqrt_above_1024 [0:2032] = '{
        0, 32, 45, 55, 64, 72, 78, 85, 91, 96, 101, 106, 111, 115, 120, 124, 128, 132, 136, 139, 143, 147, 150, 153, 157, 160, 163, 166, 169, 172, 175, 178, 181, 184, 187, 189, 192, 195, 197, 200, 202, 205, 207, 210, 212, 215, 217, 219, 222, 224, 226, 229, 231, 233, 235, 237, 239, 242, 244, 246, 248, 250, 252, 254, 256, 258, 260, 262, 264, 266, 268, 270, 272, 273, 275, 277, 279, 281, 283, 284, 286, 288, 290, 292, 293, 295, 297, 298, 300, 302, 304, 305, 307, 309, 310, 312, 314, 315, 317, 318, 320, 322, 323, 325, 326, 328, 329, 331, 333, 334, 336, 337, 339, 340, 342, 343, 345, 346, 348, 349, 351, 352, 353, 355, 356, 358, 359, 361, 362, 363, 365, 366, 368, 369, 370, 372, 373, 375, 376, 377, 379, 380, 381, 383, 384, 385, 387, 388, 389, 391, 392, 393, 395, 396, 397, 398, 400, 401, 402, 404, 405, 406, 407, 409, 410, 411, 412, 414, 415, 416, 417, 418, 420, 421, 422, 423, 425, 426, 427, 428, 429, 431, 432, 433, 434, 435, 436, 438, 439, 440, 441, 442, 443, 445, 446, 447, 448, 449, 450, 451, 453, 454, 455, 456, 457, 458, 459, 460, 462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510, 511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 532, 533, 534, 535, 535, 536, 537, 538, 539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 563, 564, 565, 566, 567, 568, 569, 570, 571, 572, 572, 573, 574, 575, 576, 577, 578, 579, 580, 580, 581, 582, 583, 584, 585, 586, 587, 587, 588, 589, 590, 591, 592, 593, 594, 594, 595, 596, 597, 598, 599, 600, 600, 601, 602, 603, 604, 605, 605, 606, 607, 608, 609, 610, 611, 611, 612, 613, 614, 615, 616, 616, 617, 618, 619, 620, 621, 621, 622, 623, 624, 625, 625, 626, 627, 628, 629, 630, 630, 631, 632, 633, 634, 634, 635, 636, 637, 638, 638, 639, 640, 641, 642, 642, 643, 644, 645, 646, 646, 647, 648, 649, 650, 650, 651, 652, 653, 653, 654, 655, 656, 657, 657, 658, 659, 660, 660, 661, 662, 663, 664, 664, 665, 666, 667, 667, 668, 669, 670, 670, 671, 672, 673, 674, 674, 675, 676, 677, 677, 678, 679, 680, 680, 681, 682, 683, 683, 684, 685, 686, 686, 687, 688, 689, 689, 690, 691, 692, 692, 693, 694, 694, 695, 696, 697, 697, 698, 699, 700, 700, 701, 702, 703, 703, 704, 705, 705, 706, 707, 708, 708, 709, 710, 711, 711, 712, 713, 713, 714, 715, 716, 716, 717, 718, 718, 719, 720, 721, 721, 722, 723, 723, 724, 725, 725, 726, 727, 728, 728, 729, 730, 730, 731, 732, 733, 733, 734, 735, 735, 736, 737, 737, 738, 739, 739, 740, 741, 742, 742, 743, 744, 744, 745, 746, 746, 747, 748, 748, 749, 750, 750, 751, 752, 753, 753, 754, 755, 755, 756, 757, 757, 758, 759, 759, 760, 761, 761, 762, 763, 763, 764, 765, 765, 766, 767, 767, 768, 769, 769, 770, 771, 771, 772, 773, 773, 774, 775, 775, 776, 777, 777, 778, 779, 779, 780, 781, 781, 782, 783, 783, 784, 784, 785, 786, 786, 787, 788, 788, 789, 790, 790, 791, 792, 792, 793, 794, 794, 795, 796, 796, 797, 797, 798, 799, 799, 800, 801, 801, 802, 803, 803, 804, 804, 805, 806, 806, 807, 808, 808, 809, 810, 810, 811, 811, 812, 813, 813, 814, 815, 815, 816, 816, 817, 818, 818, 819, 820, 820, 821, 821, 822, 823, 823, 824, 825, 825, 826, 826, 827, 828, 828, 829, 830, 830, 831, 831, 832, 833, 833, 834, 834, 835, 836, 836, 837, 838, 838, 839, 839, 840, 841, 841, 842, 842, 843, 844, 844, 845, 845, 846, 847, 847, 848, 848, 849, 850, 850, 851, 851, 852, 853, 853, 854, 854, 855, 856, 856, 857, 857, 858, 859, 859, 860, 860, 861, 862, 862, 863, 863, 864, 865, 865, 866, 866, 867, 868, 868, 869, 869, 870, 870, 871, 872, 872, 873, 873, 874, 875, 875, 876, 876, 877, 878, 878, 879, 879, 880, 880, 881, 882, 882, 883, 883, 884, 884, 885, 886, 886, 887, 887, 888, 889, 889, 890, 890, 891, 891, 892, 893, 893, 894, 894, 895, 895, 896, 897, 897, 898, 898, 899, 899, 900, 901, 901, 902, 902, 903, 903, 904, 905, 905, 906, 906, 907, 907, 908, 908, 909, 910, 910, 911, 911, 912, 912, 913, 914, 914, 915, 915, 916, 916, 917, 917, 918, 919, 919, 920, 920, 921, 921, 922, 922, 923, 924, 924, 925, 925, 926, 926, 927, 927, 928, 929, 929, 930, 930, 931, 931, 932, 932, 933, 934, 934, 935, 935, 936, 936, 937, 937, 938, 938, 939, 940, 940, 941, 941, 942, 942, 943, 943, 944, 944, 945, 945, 946, 947, 947, 948, 948, 949, 949, 950, 950, 951, 951, 952, 953, 953, 954, 954, 955, 955, 956, 956, 957, 957, 958, 958, 959, 959, 960, 961, 961, 962, 962, 963, 963, 964, 964, 965, 965, 966, 966, 967, 967, 968, 968, 969, 970, 970, 971, 971, 972, 972, 973, 973, 974, 974, 975, 975, 976, 976, 977, 977, 978, 978, 979, 980, 980, 981, 981, 982, 982, 983, 983, 984, 984, 985, 985, 986, 986, 987, 987, 988, 988, 989, 989, 990, 990, 991, 991, 992, 993, 993, 994, 994, 995, 995, 996, 996, 997, 997, 998, 998, 999, 999, 1000, 1000, 1001, 1001, 1002, 1002, 1003, 1003, 1004, 1004, 1005, 1005, 1006, 1006, 1007, 1007, 1008, 1008, 1009, 1009, 1010, 1010, 1011, 1011, 1012, 1012, 1013, 1013, 1014, 1014, 1015, 1015, 1016, 1016, 1017, 1017, 1018, 1018, 1019, 1019, 1020, 1020, 1021, 1021, 1022, 1022, 1023, 1023, 1024, 1024, 1025, 1025, 1026, 1026, 1027, 1027, 1028, 1028, 1029, 1029, 1030, 1030, 1031, 1031, 1032, 1032, 1033, 1033, 1034, 1034, 1035, 1035, 1036, 1036, 1037, 1037, 1038, 1038, 1039, 1039, 1040, 1040, 1041, 1041, 1042, 1042, 1043, 1043, 1044, 1044, 1045, 1045, 1046, 1046, 1047, 1047, 1048, 1048, 1049, 1049, 1050, 1050, 1051, 1051, 1052, 1052, 1053, 1053, 1054, 1054, 1055, 1055, 1056, 1056, 1056, 1057, 1057, 1058, 1058, 1059, 1059, 1060, 1060, 1061, 1061, 1062, 1062, 1063, 1063, 1064, 1064, 1065, 1065, 1066, 1066, 1067, 1067, 1068, 1068, 1069, 1069, 1069, 1070, 1070, 1071, 1071, 1072, 1072, 1073, 1073, 1074, 1074, 1075, 1075, 1076, 1076, 1077, 1077, 1078, 1078, 1079, 1079, 1079, 1080, 1080, 1081, 1081, 1082, 1082, 1083, 1083, 1084, 1084, 1085, 1085, 1086, 1086, 1087, 1087, 1088, 1088, 1088, 1089, 1089, 1090, 1090, 1091, 1091, 1092, 1092, 1093, 1093, 1094, 1094, 1095, 1095, 1096, 1096, 1096, 1097, 1097, 1098, 1098, 1099, 1099, 1100, 1100, 1101, 1101, 1102, 1102, 1102, 1103, 1103, 1104, 1104, 1105, 1105, 1106, 1106, 1107, 1107, 1108, 1108, 1109, 1109, 1109, 1110, 1110, 1111, 1111, 1112, 1112, 1113, 1113, 1114, 1114, 1115, 1115, 1115, 1116, 1116, 1117, 1117, 1118, 1118, 1119, 1119, 1120, 1120, 1120, 1121, 1121, 1122, 1122, 1123, 1123, 1124, 1124, 1125, 1125, 1125, 1126, 1126, 1127, 1127, 1128, 1128, 1129, 1129, 1130, 1130, 1130, 1131, 1131, 1132, 1132, 1133, 1133, 1134, 1134, 1135, 1135, 1135, 1136, 1136, 1137, 1137, 1138, 1138, 1139, 1139, 1139, 1140, 1140, 1141, 1141, 1142, 1142, 1143, 1143, 1144, 1144, 1144, 1145, 1145, 1146, 1146, 1147, 1147, 1148, 1148, 1148, 1149, 1149, 1150, 1150, 1151, 1151, 1152, 1152, 1152, 1153, 1153, 1154, 1154, 1155, 1155, 1156, 1156, 1156, 1157, 1157, 1158, 1158, 1159, 1159, 1160, 1160, 1160, 1161, 1161, 1162, 1162, 1163, 1163, 1163, 1164, 1164, 1165, 1165, 1166, 1166, 1167, 1167, 1167, 1168, 1168, 1169, 1169, 1170, 1170, 1171, 1171, 1171, 1172, 1172, 1173, 1173, 1174, 1174, 1174, 1175, 1175, 1176, 1176, 1177, 1177, 1177, 1178, 1178, 1179, 1179, 1180, 1180, 1181, 1181, 1181, 1182, 1182, 1183, 1183, 1184, 1184, 1184, 1185, 1185, 1186, 1186, 1187, 1187, 1187, 1188, 1188, 1189, 1189, 1190, 1190, 1190, 1191, 1191, 1192, 1192, 1193, 1193, 1193, 1194, 1194, 1195, 1195, 1196, 1196, 1196, 1197, 1197, 1198, 1198, 1199, 1199, 1199, 1200, 1200, 1201, 1201, 1202, 1202, 1202, 1203, 1203, 1204, 1204, 1205, 1205, 1205, 1206, 1206, 1207, 1207, 1208, 1208, 1208, 1209, 1209, 1210, 1210, 1211, 1211, 1211, 1212, 1212, 1213, 1213, 1213, 1214, 1214, 1215, 1215, 1216, 1216, 1216, 1217, 1217, 1218, 1218, 1219, 1219, 1219, 1220, 1220, 1221, 1221, 1221, 1222, 1222, 1223, 1223, 1224, 1224, 1224, 1225, 1225, 1226, 1226, 1226, 1227, 1227, 1228, 1228, 1229, 1229, 1229, 1230, 1230, 1231, 1231, 1231, 1232, 1232, 1233, 1233, 1234, 1234, 1234, 1235, 1235, 1236, 1236, 1236, 1237, 1237, 1238, 1238, 1239, 1239, 1239, 1240, 1240, 1241, 1241, 1241, 1242, 1242, 1243, 1243, 1243, 1244, 1244, 1245, 1245, 1246, 1246, 1246, 1247, 1247, 1248, 1248, 1248, 1249, 1249, 1250, 1250, 1250, 1251, 1251, 1252, 1252, 1253, 1253, 1253, 1254, 1254, 1255, 1255, 1255, 1256, 1256, 1257, 1257, 1257, 1258, 1258, 1259, 1259, 1259, 1260, 1260, 1261, 1261, 1261, 1262, 1262, 1263, 1263, 1263, 1264, 1264, 1265, 1265, 1266, 1266, 1266, 1267, 1267, 1268, 1268, 1268, 1269, 1269, 1270, 1270, 1270, 1271, 1271, 1272, 1272, 1272, 1273, 1273, 1274, 1274, 1274, 1275, 1275, 1276, 1276, 1276, 1277, 1277, 1278, 1278, 1278, 1279, 1279, 1280, 1280, 1280, 1281, 1281, 1282, 1282, 1282, 1283, 1283, 1284, 1284, 1284, 1285, 1285, 1286, 1286, 1286, 1287, 1287, 1288, 1288, 1288, 1289, 1289, 1290, 1290, 1290, 1291, 1291, 1292, 1292, 1292, 1293, 1293, 1294, 1294, 1294, 1295, 1295, 1296, 1296, 1296, 1297, 1297, 1297, 1298, 1298, 1299, 1299, 1299, 1300, 1300, 1301, 1301, 1301, 1302, 1302, 1303, 1303, 1303, 1304, 1304, 1305, 1305, 1305, 1306, 1306, 1307, 1307, 1307, 1308, 1308, 1308, 1309, 1309, 1310, 1310, 1310, 1311, 1311, 1312, 1312, 1312, 1313, 1313, 1314, 1314, 1314, 1315, 1315, 1316, 1316, 1316, 1317, 1317, 1317, 1318, 1318, 1319, 1319, 1319, 1320, 1320, 1321, 1321, 1321, 1322, 1322, 1322, 1323, 1323, 1324, 1324, 1324, 1325, 1325, 1326, 1326, 1326, 1327, 1327, 1328, 1328, 1328, 1329, 1329, 1329, 1330, 1330, 1331, 1331, 1331, 1332, 1332, 1333, 1333, 1333, 1334, 1334, 1334, 1335, 1335, 1336, 1336, 1336, 1337, 1337, 1338, 1338, 1338, 1339, 1339, 1339, 1340, 1340, 1341, 1341, 1341, 1342, 1342, 1342, 1343, 1343, 1344, 1344, 1344, 1345, 1345, 1346, 1346, 1346, 1347, 1347, 1347, 1348, 1348, 1349, 1349, 1349, 1350, 1350, 1350, 1351, 1351, 1352, 1352, 1352, 1353, 1353, 1353, 1354, 1354, 1355, 1355, 1355, 1356, 1356, 1357, 1357, 1357, 1358, 1358, 1358, 1359, 1359, 1360, 1360, 1360, 1361, 1361, 1361, 1362, 1362, 1363, 1363, 1363, 1364, 1364, 1364, 1365, 1365, 1366, 1366, 1366, 1367, 1367, 1367, 1368, 1368, 1369, 1369, 1369, 1370, 1370, 1370, 1371, 1371, 1372, 1372, 1372, 1373, 1373, 1373, 1374, 1374, 1375, 1375, 1375, 1376, 1376, 1376, 1377, 1377, 1377, 1378, 1378, 1379, 1379, 1379, 1380, 1380, 1380, 1381, 1381, 1382, 1382, 1382, 1383, 1383, 1383, 1384, 1384, 1385, 1385, 1385, 1386, 1386, 1386, 1387, 1387, 1387, 1388, 1388, 1389, 1389, 1389, 1390, 1390, 1390, 1391, 1391, 1392, 1392, 1392, 1393, 1393, 1393, 1394, 1394, 1394, 1395, 1395, 1396, 1396, 1396, 1397, 1397, 1397, 1398, 1398, 1399, 1399, 1399, 1400, 1400, 1400, 1401, 1401, 1401, 1402, 1402, 1403, 1403, 1403, 1404, 1404, 1404, 1405, 1405, 1405, 1406, 1406, 1407, 1407, 1407, 1408, 1408, 1408, 1409, 1409, 1409, 1410, 1410, 1411, 1411, 1411, 1412, 1412, 1412, 1413, 1413, 1413, 1414, 1414, 1415, 1415, 1415, 1416, 1416, 1416, 1417, 1417, 1417, 1418, 1418, 1419, 1419, 1419, 1420, 1420, 1420, 1421, 1421, 1421, 1422, 1422, 1422, 1423, 1423, 1424, 1424, 1424, 1425, 1425, 1425, 1426, 1426, 1426, 1427, 1427, 1428, 1428, 1428, 1429, 1429, 1429, 1430, 1430, 1430, 1431, 1431, 1431, 1432, 1432, 1433, 1433, 1433, 1434, 1434, 1434, 1435, 1435, 1435, 1436, 1436, 1436, 1437, 1437, 1438, 1438, 1438, 1439, 1439, 1439, 1440, 1440, 1440, 1441, 1441, 1441, 1442, 1442, 1442 
    };

    logic [10:0] index;
    logic [9:0]  offset;
    logic [10:0] base, next;
    logic [20:0] adjustment;

    always_comb begin
        index   = 0;
        offset  = 0;
        base    = 0;
        next    = 0;
        adjustment = 0;
        
        if (value < 1024) begin
            sqrt = sqrt_below_1024[value];
        end
        else begin
            index  = value >> 10;
            offset = value[9:0];

            base = sqrt_above_1024[index];
            next = (index < 2032)? sqrt_above_1024[index + 1] : base;
            
            adjustment = ((next - base) * offset) >> 10;
            sqrt = base + adjustment;
        end
    end

endmodule
